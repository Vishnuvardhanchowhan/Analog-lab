zener regulator
.subckt ZENER_12 1 2
d1 1 2 df
dz 3 1 dr
vz 2 3 10.8
.model df D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n)
.model dr D ( IS=5.49f RS=50 N=1.77 )
.ends
r1  1 2 470
vs 2 3 0
x1 4 3 ZENER_12
vze 4 0 0
r2 3 5 500
vl 5 0 0
vin 1 0
.dc vin 15 25 0.5
.control
run
print v(3)
plot v(3)
.endc
.end


