instrumentation amplifier
.subckt ua741    1  2  3  4  5
c1   11 12 8.661E-12
c2    6  7 30.00E-12
dc    5 53 dx
de   54  5 dx
dlp  90 91 dx
dln  92 90 dx
dp    4  3 dx
egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
ga    6  0 11 12 188.5E-6
gcm   0  6 10 99 5.961E-9
iee  10  4 dc 15.16E-6
hlim 90  0 vlim 1K
q1   11  2 13 qx
q2   12  1 14 qx
r2    6  9 100.0E3
rc1   3 11 5.305E3
rc2   3 12 5.305E3
re1  13 10 1.836E3
re2  14 10 1.836E3
ree  10 99 13.19E6
ro1   8  5 50
ro2   7 99 100
rp    3  4 18.16E3
vb    9  0 dc 0
vc    3 53 dc 1
ve   54  4 dc 1
vlim  7  8 dc 0
vlp  91  0 dc 40
vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
vcm 1 0 dc 
vi1 1 2 0
vi2 1 4 0
x3 2 3 6 7 8 ua741
x2 4 5 9 10 11 ua741
r10 3 5 2.21k
r5 5 11 10k
vcc31 6 0 15v
vcc32 7 0 -15v
vcc21 9 0 15v
vcc22 10 0 -15v
r6 3 8 10k
r1 8 12 10k
r2 12 13 10k
r3 11 14 10k
r4 14 15 10k
vref 15 0 0
x1 14 12 16 17 13 ua741
vcc11 16 0 15v
vcc12 17 0 -15v
.dc vcm -2 2 1m
.control
run
plot v(13)
.endc
.end 
