schmitt trigger circuit
.subckt ua741    1  2  3  4  5
c1   11 12 8.661E-12
c2    6  7 30.00E-12
dc    5 53 dx
de   54  5 dx
dlp  90 91 dx
dln  92 90 dx
dp    4  3 dx
egnd 99  0 poly(2) (3,0) (4,0) 0 .5 .5
fb    7 99 poly(5) vb vc ve vlp vln 0 10.61E6 -10E6 10E6 10E6 -10E6
ga    6  0 11 12 188.5E-6
gcm   0  6 10 99 5.961E-9
iee  10  4 dc 15.16E-6
hlim 90  0 vlim 1K
q1   11  2 13 qx
q2   12  1 14 qx
r2    6  9 100.0E3
rc1   3 11 5.305E3
rc2   3 12 5.305E3
re1  13 10 1.836E3
re2  14 10 1.836E3
ree  10 99 13.19E6
ro1   8  5 50
ro2   7 99 100
rp    3  4 18.16E3
vb    9  0 dc 0
vc    3 53 dc 1
ve   54  4 dc 1
vlim  7  8 dc 0
vlp  91  0 dc 40
vln   0 92 dc 40
.model dx D(Is=800.0E-18 Rs=1)
.model qx NPN(Is=800.0E-18 Bf=93.75)
.ends
.subckt ZENER_12 1 2
d1 1 2 df
dz 3 1 dr
vz 2 3 3.5
.model df D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n)
.model dr D ( IS=5.49f RS=50 N=1.77 )
.ends

vin 1 0 sin(0 6 1k 0 0)
x1 5 1 6 7 2 ua741
ro 2 3 1k
r2 3 5 10k
r1 5 8 10k
va 8 0 -3v
x2 3 4 ZENER_12
x3 0 4 ZENER_12
vdd1 6 0 15v
vdd2 7 0 -15v
.tran 0.01u 4m
.control
run 
plot v(3) v(1)
.endc 
.end

